(*blackbox*)
module OTA_2stage_macro (
`ifdef USE_POWER_PINS
    inout VDD,
    inout VSS,
`endif
);
endmodule // OTA_2stage
